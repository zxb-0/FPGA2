library verilog;
use verilog.vl_types.all;
entity final_top_tb is
end final_top_tb;
